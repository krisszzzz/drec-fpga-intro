
`define CBU_OP_EQ 3'b000
`define CBU_OP_NE 3'b001
`define CBU_OP_LT 3'b010
`define CBU_OP_GE 3'b011
`define CBU_OP_LTU 3'b100
`define CBU_OP_GEU 3'b101
`define CBU_OP_INV 3'b111